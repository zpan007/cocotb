package test_pkg;

    typedef struct packed {
        logic                           status0;
        logic                           status1;
        logic                           status2;
    } test_status_t;



endpackage: test_pkg
